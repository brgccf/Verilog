module hello;
	initial begin
		$display ("Hello World!");
		$display ("Hello World!");
		#10 $finish;
	end

endmodule